Bit #(12) csr_addr_vstart = 12'h008;
Bit #(12) csr_addr_vxsat  = 12'h009;
Bit #(12) csr_addr_vxrm   = 12'h000A;
Bit #(12) csr_addr_vl     = 12'hC20;
Bit #(12) csr_addr_vtype  = 12'hC21;
Bit #(12) csr_addr_vlenb  = 12'hC22;